LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY wav_rom IS
PORT (
      CLOCK          : IN  STD_LOGIC;
      ADDR_R         : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
      DATA_OUT       : OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
      );
END wav_rom;

ARCHITECTURE Behavioral OF wav_rom IS

  TYPE rom_type IS ARRAY (0 TO 44099) OF SIGNED (10 DOWNTO 0);
  SIGNAL memory : rom_type := (
    TO_SIGNED(   0, 11), TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED( 657, 11), TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED( 549, 11), TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11), TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11), TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11), TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED( 381, 11), TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED( 718, 11), TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED( 218, 11), TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11), TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11), TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED( -20, 11), TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED( 648, 11), TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED( 562, 11), TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11), TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11), TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11), TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED( 364, 11), TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED( 720, 11), TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED( 237, 11), TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11), TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11), TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED( -41, 11), TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED( 639, 11), TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED( 575, 11), TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11), TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),
    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),
    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),
    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),
    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),
    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),
    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),
    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),
    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),
    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),
    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),
    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),
    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),
    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),
    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),
    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),
    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),
    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),
    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),
    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),
    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),
    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),
    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),
    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),
    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),
    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),
    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),
    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),
    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),
    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),
    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),
    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),
    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),
    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),
    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),
    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),
    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),
    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),
    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),
    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),
    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),
    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),
    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),
    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),
    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),
    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),
    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),
    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),
    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),
    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),
    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),
    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),
    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),
    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),
    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),
    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),
    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),
    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),
    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),
    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),
    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),
    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),
    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),
    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),
    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),
    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),
    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),
    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),
    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),
    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),
    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),
    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),
    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),
    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),
    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),
    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),
    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),
    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),
    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),
    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),
    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),
    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),
    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),
    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),
    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),
    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),
    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),
    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),
    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),
    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),
    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),
    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),
    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),
    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),
    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),
    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),
    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),
    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),
    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),
    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),
    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),
    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),
    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),
    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),
    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),
    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),
    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),
    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),
    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),
    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),
    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),
    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),
    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),
    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),
    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),
    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),
    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),
    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),
    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),
    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),
    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),
    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),
    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),
    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),
    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),
    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),
    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),
    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),
    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),
    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),
    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),
    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),
    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),
    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),
    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),
    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),
    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),
    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),
    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),
    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),
    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),
    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),
    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),
    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),
    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),
    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),
    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),
    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),
    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),
    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),
    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),
    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),
    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),
    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),
    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),
    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),
    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),
    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),
    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),
    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),
    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),
    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),
    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),
    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),
    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),
    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),
    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),
    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),
    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),
    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),
    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),
    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),
    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),
    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),
    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),
    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),
    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),
    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),
    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),
    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),
    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),
    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),
    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),
    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),
    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),
    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),
    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),
    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),
    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),
    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),
    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),
    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),
    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),
    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),
    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),
    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),
    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),
    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),
    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),
    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),
    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),
    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),
    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),
    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),
    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),
    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),
    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),
    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),
    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),
    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),
    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),
    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),
    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),
    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),
    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),
    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),
    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),
    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),
    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),
    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),
    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),
    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),
    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),
    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),
    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),
    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),
    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),
    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),
    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),
    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),
    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),
    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),
    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),
    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),
    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),
    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),
    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),
    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),
    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),
    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),
    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),
    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),
    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),
    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),
    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),
    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),
    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),
    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),
    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),
    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),
    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),
    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),
    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),
    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),
    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),
    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),
    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),
    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),
    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),
    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),
    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),
    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),
    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),
    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),
    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),
    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),
    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),
    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),
    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),
    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),
    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),
    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),
    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),
    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),
    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),    TO_SIGNED(546, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),    TO_SIGNED(660, 11),
    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),    TO_SIGNED(5, 11),
    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),    TO_SIGNED(-655, 11),
    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),    TO_SIGNED(-553, 11),
    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),    TO_SIGNED(193, 11),
    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),    TO_SIGNED(714, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),    TO_SIGNED(403, 11),
    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),    TO_SIGNED(-377, 11),
    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),    TO_SIGNED(-223, 11),
    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),    TO_SIGNED(532, 11),
    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),    TO_SIGNED(668, 11),
    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),    TO_SIGNED(25, 11),
    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),    TO_SIGNED(-646, 11),
    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),    TO_SIGNED(-566, 11),
    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),    TO_SIGNED(173, 11),
    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),    TO_SIGNED(711, 11),
    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),    TO_SIGNED(420, 11),
    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-359, 11),
    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),    TO_SIGNED(-242, 11),
    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),    TO_SIGNED(518, 11),
    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),    TO_SIGNED(675, 11),
    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),    TO_SIGNED(46, 11),
    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),    TO_SIGNED(-637, 11),
    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),    TO_SIGNED(-578, 11),
    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),    TO_SIGNED(153, 11),
    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),    TO_SIGNED(707, 11),
    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),    TO_SIGNED(437, 11),
    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),    TO_SIGNED(-341, 11),
    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),    TO_SIGNED(-722, 11),
    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),    TO_SIGNED(-262, 11),
    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),    TO_SIGNED(503, 11),
    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),    TO_SIGNED(683, 11),
    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),    TO_SIGNED(66, 11),
    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),    TO_SIGNED(-627, 11),
    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),    TO_SIGNED(133, 11),
    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),    TO_SIGNED(702, 11),
    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),    TO_SIGNED(453, 11),
    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),    TO_SIGNED(-323, 11),
    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-281, 11),
    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),    TO_SIGNED(488, 11),
    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),    TO_SIGNED(689, 11),
    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),    TO_SIGNED(87, 11),
    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),    TO_SIGNED(-616, 11),
    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),    TO_SIGNED(-602, 11),
    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),    TO_SIGNED(113, 11),
    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),    TO_SIGNED(469, 11),
    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),    TO_SIGNED(-304, 11),
    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-724, 11),
    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),    TO_SIGNED(-300, 11),
    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(203, 11),    TO_SIGNED(300, 11),    TO_SIGNED(390, 11),    TO_SIGNED(473, 11),
    TO_SIGNED(546, 11),    TO_SIGNED(608, 11),    TO_SIGNED(657, 11),    TO_SIGNED(694, 11),    TO_SIGNED(716, 11),    TO_SIGNED(724, 11),    TO_SIGNED(717, 11),    TO_SIGNED(695, 11),
    TO_SIGNED(660, 11),    TO_SIGNED(611, 11),    TO_SIGNED(549, 11),    TO_SIGNED(477, 11),    TO_SIGNED(395, 11),    TO_SIGNED(304, 11),    TO_SIGNED(208, 11),    TO_SIGNED(107, 11),
    TO_SIGNED(5, 11),    TO_SIGNED(-97, 11),    TO_SIGNED(-198, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-386, 11),    TO_SIGNED(-469, 11),    TO_SIGNED(-542, 11),    TO_SIGNED(-605, 11),
    TO_SIGNED(-655, 11),    TO_SIGNED(-692, 11),    TO_SIGNED(-715, 11),    TO_SIGNED(-724, 11),    TO_SIGNED(-717, 11),    TO_SIGNED(-697, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-613, 11),
    TO_SIGNED(-553, 11),    TO_SIGNED(-481, 11),    TO_SIGNED(-399, 11),    TO_SIGNED(-309, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-10, 11),    TO_SIGNED(92, 11),
    TO_SIGNED(193, 11),    TO_SIGNED(290, 11),    TO_SIGNED(381, 11),    TO_SIGNED(465, 11),    TO_SIGNED(539, 11),    TO_SIGNED(602, 11),    TO_SIGNED(653, 11),    TO_SIGNED(691, 11),
    TO_SIGNED(714, 11),    TO_SIGNED(723, 11),    TO_SIGNED(718, 11),    TO_SIGNED(698, 11),    TO_SIGNED(664, 11),    TO_SIGNED(616, 11),    TO_SIGNED(556, 11),    TO_SIGNED(484, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(314, 11),    TO_SIGNED(218, 11),    TO_SIGNED(118, 11),    TO_SIGNED(15, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-286, 11),
    TO_SIGNED(-377, 11),    TO_SIGNED(-461, 11),    TO_SIGNED(-536, 11),    TO_SIGNED(-599, 11),    TO_SIGNED(-651, 11),    TO_SIGNED(-689, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-719, 11),    TO_SIGNED(-699, 11),    TO_SIGNED(-666, 11),    TO_SIGNED(-619, 11),    TO_SIGNED(-559, 11),    TO_SIGNED(-488, 11),    TO_SIGNED(-407, 11),    TO_SIGNED(-318, 11),
    TO_SIGNED(-223, 11),    TO_SIGNED(-123, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(82, 11),    TO_SIGNED(183, 11),    TO_SIGNED(281, 11),    TO_SIGNED(373, 11),    TO_SIGNED(457, 11),
    TO_SIGNED(532, 11),    TO_SIGNED(596, 11),    TO_SIGNED(648, 11),    TO_SIGNED(688, 11),    TO_SIGNED(713, 11),    TO_SIGNED(723, 11),    TO_SIGNED(719, 11),    TO_SIGNED(701, 11),
    TO_SIGNED(668, 11),    TO_SIGNED(621, 11),    TO_SIGNED(562, 11),    TO_SIGNED(492, 11),    TO_SIGNED(412, 11),    TO_SIGNED(323, 11),    TO_SIGNED(228, 11),    TO_SIGNED(128, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-178, 11),    TO_SIGNED(-276, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-453, 11),    TO_SIGNED(-529, 11),    TO_SIGNED(-593, 11),
    TO_SIGNED(-646, 11),    TO_SIGNED(-686, 11),    TO_SIGNED(-712, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-702, 11),    TO_SIGNED(-670, 11),    TO_SIGNED(-624, 11),
    TO_SIGNED(-566, 11),    TO_SIGNED(-496, 11),    TO_SIGNED(-416, 11),    TO_SIGNED(-328, 11),    TO_SIGNED(-233, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-30, 11),    TO_SIGNED(72, 11),
    TO_SIGNED(173, 11),    TO_SIGNED(271, 11),    TO_SIGNED(364, 11),    TO_SIGNED(449, 11),    TO_SIGNED(525, 11),    TO_SIGNED(590, 11),    TO_SIGNED(644, 11),    TO_SIGNED(684, 11),
    TO_SIGNED(711, 11),    TO_SIGNED(723, 11),    TO_SIGNED(720, 11),    TO_SIGNED(703, 11),    TO_SIGNED(672, 11),    TO_SIGNED(627, 11),    TO_SIGNED(569, 11),    TO_SIGNED(500, 11),
    TO_SIGNED(420, 11),    TO_SIGNED(332, 11),    TO_SIGNED(237, 11),    TO_SIGNED(138, 11),    TO_SIGNED(36, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-168, 11),    TO_SIGNED(-266, 11),
    TO_SIGNED(-359, 11),    TO_SIGNED(-445, 11),    TO_SIGNED(-521, 11),    TO_SIGNED(-587, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-683, 11),    TO_SIGNED(-710, 11),    TO_SIGNED(-723, 11),
    TO_SIGNED(-721, 11),    TO_SIGNED(-704, 11),    TO_SIGNED(-674, 11),    TO_SIGNED(-629, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-503, 11),    TO_SIGNED(-424, 11),    TO_SIGNED(-337, 11),
    TO_SIGNED(-242, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(61, 11),    TO_SIGNED(163, 11),    TO_SIGNED(262, 11),    TO_SIGNED(355, 11),    TO_SIGNED(441, 11),
    TO_SIGNED(518, 11),    TO_SIGNED(584, 11),    TO_SIGNED(639, 11),    TO_SIGNED(681, 11),    TO_SIGNED(709, 11),    TO_SIGNED(722, 11),    TO_SIGNED(721, 11),    TO_SIGNED(705, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(632, 11),    TO_SIGNED(575, 11),    TO_SIGNED(507, 11),    TO_SIGNED(428, 11),    TO_SIGNED(341, 11),    TO_SIGNED(247, 11),    TO_SIGNED(148, 11),
    TO_SIGNED(46, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-257, 11),    TO_SIGNED(-350, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-514, 11),    TO_SIGNED(-581, 11),
    TO_SIGNED(-637, 11),    TO_SIGNED(-679, 11),    TO_SIGNED(-708, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-722, 11),    TO_SIGNED(-707, 11),    TO_SIGNED(-677, 11),    TO_SIGNED(-634, 11),
    TO_SIGNED(-578, 11),    TO_SIGNED(-511, 11),    TO_SIGNED(-433, 11),    TO_SIGNED(-346, 11),    TO_SIGNED(-252, 11),    TO_SIGNED(-153, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(153, 11),    TO_SIGNED(252, 11),    TO_SIGNED(346, 11),    TO_SIGNED(433, 11),    TO_SIGNED(511, 11),    TO_SIGNED(578, 11),    TO_SIGNED(634, 11),    TO_SIGNED(677, 11),
    TO_SIGNED(707, 11),    TO_SIGNED(722, 11),    TO_SIGNED(722, 11),    TO_SIGNED(708, 11),    TO_SIGNED(679, 11),    TO_SIGNED(637, 11),    TO_SIGNED(581, 11),    TO_SIGNED(514, 11),
    TO_SIGNED(437, 11),    TO_SIGNED(350, 11),    TO_SIGNED(257, 11),    TO_SIGNED(158, 11),    TO_SIGNED(56, 11),    TO_SIGNED(-46, 11),    TO_SIGNED(-148, 11),    TO_SIGNED(-247, 11),
    TO_SIGNED(-341, 11),    TO_SIGNED(-428, 11),    TO_SIGNED(-507, 11),    TO_SIGNED(-575, 11),    TO_SIGNED(-632, 11),    TO_SIGNED(-675, 11),    TO_SIGNED(-705, 11),    TO_SIGNED(-721, 11),
    TO_SIGNED(-722, 11),    TO_SIGNED(-709, 11),    TO_SIGNED(-681, 11),    TO_SIGNED(-639, 11),    TO_SIGNED(-584, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-441, 11),    TO_SIGNED(-355, 11),
    TO_SIGNED(-262, 11),    TO_SIGNED(-163, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(41, 11),    TO_SIGNED(143, 11),    TO_SIGNED(242, 11),    TO_SIGNED(337, 11),    TO_SIGNED(424, 11),
    TO_SIGNED(503, 11),    TO_SIGNED(572, 11),    TO_SIGNED(629, 11),    TO_SIGNED(674, 11),    TO_SIGNED(704, 11),    TO_SIGNED(721, 11),    TO_SIGNED(723, 11),    TO_SIGNED(710, 11),
    TO_SIGNED(683, 11),    TO_SIGNED(641, 11),    TO_SIGNED(587, 11),    TO_SIGNED(521, 11),    TO_SIGNED(445, 11),    TO_SIGNED(359, 11),    TO_SIGNED(266, 11),    TO_SIGNED(168, 11),
    TO_SIGNED(66, 11),    TO_SIGNED(-36, 11),    TO_SIGNED(-138, 11),    TO_SIGNED(-237, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-420, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-569, 11),
    TO_SIGNED(-627, 11),    TO_SIGNED(-672, 11),    TO_SIGNED(-703, 11),    TO_SIGNED(-720, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-711, 11),    TO_SIGNED(-684, 11),    TO_SIGNED(-644, 11),
    TO_SIGNED(-590, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-364, 11),    TO_SIGNED(-271, 11),    TO_SIGNED(-173, 11),    TO_SIGNED(-72, 11),    TO_SIGNED(30, 11),
    TO_SIGNED(133, 11),    TO_SIGNED(233, 11),    TO_SIGNED(328, 11),    TO_SIGNED(416, 11),    TO_SIGNED(496, 11),    TO_SIGNED(566, 11),    TO_SIGNED(624, 11),    TO_SIGNED(670, 11),
    TO_SIGNED(702, 11),    TO_SIGNED(720, 11),    TO_SIGNED(723, 11),    TO_SIGNED(712, 11),    TO_SIGNED(686, 11),    TO_SIGNED(646, 11),    TO_SIGNED(593, 11),    TO_SIGNED(529, 11),
    TO_SIGNED(453, 11),    TO_SIGNED(368, 11),    TO_SIGNED(276, 11),    TO_SIGNED(178, 11),    TO_SIGNED(77, 11),    TO_SIGNED(-25, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-228, 11),
    TO_SIGNED(-323, 11),    TO_SIGNED(-412, 11),    TO_SIGNED(-492, 11),    TO_SIGNED(-562, 11),    TO_SIGNED(-621, 11),    TO_SIGNED(-668, 11),    TO_SIGNED(-701, 11),    TO_SIGNED(-719, 11),
    TO_SIGNED(-723, 11),    TO_SIGNED(-713, 11),    TO_SIGNED(-688, 11),    TO_SIGNED(-648, 11),    TO_SIGNED(-596, 11),    TO_SIGNED(-532, 11),    TO_SIGNED(-457, 11),    TO_SIGNED(-373, 11),
    TO_SIGNED(-281, 11),    TO_SIGNED(-183, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(20, 11),    TO_SIGNED(123, 11),    TO_SIGNED(223, 11),    TO_SIGNED(318, 11),    TO_SIGNED(407, 11),
    TO_SIGNED(488, 11),    TO_SIGNED(559, 11),    TO_SIGNED(619, 11),    TO_SIGNED(666, 11),    TO_SIGNED(699, 11),    TO_SIGNED(719, 11),    TO_SIGNED(723, 11),    TO_SIGNED(713, 11),
    TO_SIGNED(689, 11),    TO_SIGNED(651, 11),    TO_SIGNED(599, 11),    TO_SIGNED(536, 11),    TO_SIGNED(461, 11),    TO_SIGNED(377, 11),    TO_SIGNED(286, 11),    TO_SIGNED(188, 11),
    TO_SIGNED(87, 11),    TO_SIGNED(-15, 11),    TO_SIGNED(-118, 11),    TO_SIGNED(-218, 11),    TO_SIGNED(-314, 11),    TO_SIGNED(-403, 11),    TO_SIGNED(-484, 11),    TO_SIGNED(-556, 11),
    TO_SIGNED(-616, 11),    TO_SIGNED(-664, 11),    TO_SIGNED(-698, 11),    TO_SIGNED(-718, 11),    TO_SIGNED(-723, 11),    TO_SIGNED(-714, 11),    TO_SIGNED(-691, 11),    TO_SIGNED(-653, 11),
    TO_SIGNED(-602, 11),    TO_SIGNED(-539, 11),    TO_SIGNED(-465, 11),    TO_SIGNED(-381, 11),    TO_SIGNED(-290, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(10, 11),
    TO_SIGNED(113, 11),    TO_SIGNED(213, 11),    TO_SIGNED(309, 11),    TO_SIGNED(399, 11),    TO_SIGNED(481, 11),    TO_SIGNED(553, 11),    TO_SIGNED(613, 11),    TO_SIGNED(662, 11),
    TO_SIGNED(697, 11),    TO_SIGNED(717, 11),    TO_SIGNED(724, 11),    TO_SIGNED(715, 11),    TO_SIGNED(692, 11),    TO_SIGNED(655, 11),    TO_SIGNED(605, 11),    TO_SIGNED(542, 11),
    TO_SIGNED(469, 11),    TO_SIGNED(386, 11),    TO_SIGNED(295, 11),    TO_SIGNED(198, 11),    TO_SIGNED(97, 11),    TO_SIGNED(-5, 11),    TO_SIGNED(-107, 11),    TO_SIGNED(-208, 11),
    TO_SIGNED(-304, 11),    TO_SIGNED(-395, 11),    TO_SIGNED(-477, 11),    TO_SIGNED(-549, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-660, 11),    TO_SIGNED(-695, 11),    TO_SIGNED(-717, 11),
    TO_SIGNED(-724, 11),    TO_SIGNED(-716, 11),    TO_SIGNED(-694, 11),    TO_SIGNED(-657, 11),    TO_SIGNED(-608, 11),    TO_SIGNED(-546, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-390, 11),
    TO_SIGNED(-300, 11),    TO_SIGNED(-203, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(0, 11),    TO_SIGNED(102, 11),    TO_SIGNED(202, 11),    TO_SIGNED(298, 11),    TO_SIGNED(387, 11),
    TO_SIGNED(467, 11),    TO_SIGNED(538, 11),    TO_SIGNED(598, 11),    TO_SIGNED(645, 11),    TO_SIGNED(680, 11),    TO_SIGNED(700, 11),    TO_SIGNED(706, 11),    TO_SIGNED(697, 11),
    TO_SIGNED(675, 11),    TO_SIGNED(639, 11),    TO_SIGNED(590, 11),    TO_SIGNED(529, 11),    TO_SIGNED(458, 11),    TO_SIGNED(378, 11),    TO_SIGNED(291, 11),    TO_SIGNED(199, 11),
    TO_SIGNED(102, 11),    TO_SIGNED(4, 11),    TO_SIGNED(-92, 11),    TO_SIGNED(-187, 11),    TO_SIGNED(-278, 11),    TO_SIGNED(-363, 11),    TO_SIGNED(-440, 11),    TO_SIGNED(-508, 11),
    TO_SIGNED(-565, 11),    TO_SIGNED(-611, 11),    TO_SIGNED(-643, 11),    TO_SIGNED(-663, 11),    TO_SIGNED(-669, 11),    TO_SIGNED(-662, 11),    TO_SIGNED(-641, 11),    TO_SIGNED(-608, 11),
    TO_SIGNED(-562, 11),    TO_SIGNED(-505, 11),    TO_SIGNED(-438, 11),    TO_SIGNED(-363, 11),    TO_SIGNED(-280, 11),    TO_SIGNED(-193, 11),    TO_SIGNED(-102, 11),    TO_SIGNED(-9, 11),
    TO_SIGNED(83, 11),    TO_SIGNED(173, 11),    TO_SIGNED(259, 11),    TO_SIGNED(340, 11),    TO_SIGNED(413, 11),    TO_SIGNED(478, 11),    TO_SIGNED(532, 11),    TO_SIGNED(576, 11),
    TO_SIGNED(608, 11),    TO_SIGNED(627, 11),    TO_SIGNED(633, 11),    TO_SIGNED(627, 11),    TO_SIGNED(608, 11),    TO_SIGNED(576, 11),    TO_SIGNED(534, 11),    TO_SIGNED(480, 11),
    TO_SIGNED(417, 11),    TO_SIGNED(346, 11),    TO_SIGNED(269, 11),    TO_SIGNED(186, 11),    TO_SIGNED(100, 11),    TO_SIGNED(13, 11),    TO_SIGNED(-74, 11),    TO_SIGNED(-159, 11),
    TO_SIGNED(-241, 11),    TO_SIGNED(-317, 11),    TO_SIGNED(-387, 11),    TO_SIGNED(-448, 11),    TO_SIGNED(-500, 11),    TO_SIGNED(-541, 11),    TO_SIGNED(-572, 11),    TO_SIGNED(-590, 11),
    TO_SIGNED(-597, 11),    TO_SIGNED(-591, 11),    TO_SIGNED(-574, 11),    TO_SIGNED(-545, 11),    TO_SIGNED(-505, 11),    TO_SIGNED(-455, 11),    TO_SIGNED(-396, 11),    TO_SIGNED(-330, 11),
    TO_SIGNED(-257, 11),    TO_SIGNED(-179, 11),    TO_SIGNED(-98, 11),    TO_SIGNED(-16, 11),    TO_SIGNED(65, 11),    TO_SIGNED(146, 11),    TO_SIGNED(223, 11),    TO_SIGNED(295, 11),
    TO_SIGNED(361, 11),    TO_SIGNED(419, 11),    TO_SIGNED(468, 11),    TO_SIGNED(507, 11),    TO_SIGNED(536, 11),    TO_SIGNED(554, 11),    TO_SIGNED(561, 11),    TO_SIGNED(556, 11),
    TO_SIGNED(540, 11),    TO_SIGNED(513, 11),    TO_SIGNED(476, 11),    TO_SIGNED(430, 11),    TO_SIGNED(375, 11),    TO_SIGNED(313, 11),    TO_SIGNED(244, 11),    TO_SIGNED(172, 11),
    TO_SIGNED(96, 11),    TO_SIGNED(19, 11),    TO_SIGNED(-57, 11),    TO_SIGNED(-133, 11),    TO_SIGNED(-205, 11),    TO_SIGNED(-273, 11),    TO_SIGNED(-335, 11),    TO_SIGNED(-389, 11),
    TO_SIGNED(-436, 11),    TO_SIGNED(-473, 11),    TO_SIGNED(-501, 11),    TO_SIGNED(-518, 11),    TO_SIGNED(-525, 11),    TO_SIGNED(-520, 11),    TO_SIGNED(-506, 11),    TO_SIGNED(-481, 11),
    TO_SIGNED(-447, 11),    TO_SIGNED(-404, 11),    TO_SIGNED(-353, 11),    TO_SIGNED(-295, 11),    TO_SIGNED(-232, 11),    TO_SIGNED(-164, 11),    TO_SIGNED(-93, 11),    TO_SIGNED(-21, 11),
    TO_SIGNED(50, 11),    TO_SIGNED(120, 11),    TO_SIGNED(188, 11),    TO_SIGNED(251, 11),    TO_SIGNED(309, 11),    TO_SIGNED(361, 11),    TO_SIGNED(404, 11),    TO_SIGNED(439, 11),
    TO_SIGNED(465, 11),    TO_SIGNED(482, 11),    TO_SIGNED(488, 11),    TO_SIGNED(485, 11),    TO_SIGNED(472, 11),    TO_SIGNED(449, 11),    TO_SIGNED(418, 11),    TO_SIGNED(378, 11),
    TO_SIGNED(331, 11),    TO_SIGNED(277, 11),    TO_SIGNED(218, 11),    TO_SIGNED(155, 11),    TO_SIGNED(90, 11),    TO_SIGNED(23, 11),    TO_SIGNED(-43, 11),    TO_SIGNED(-109, 11),
    TO_SIGNED(-171, 11),    TO_SIGNED(-230, 11),    TO_SIGNED(-284, 11),    TO_SIGNED(-332, 11),    TO_SIGNED(-373, 11),    TO_SIGNED(-406, 11),    TO_SIGNED(-430, 11),    TO_SIGNED(-446, 11),
    TO_SIGNED(-452, 11),    TO_SIGNED(-449, 11),    TO_SIGNED(-437, 11),    TO_SIGNED(-417, 11),    TO_SIGNED(-388, 11),    TO_SIGNED(-351, 11),    TO_SIGNED(-308, 11),    TO_SIGNED(-259, 11),
    TO_SIGNED(-204, 11),    TO_SIGNED(-147, 11),    TO_SIGNED(-86, 11),    TO_SIGNED(-24, 11),    TO_SIGNED(37, 11),    TO_SIGNED(97, 11),    TO_SIGNED(155, 11),    TO_SIGNED(210, 11),
    TO_SIGNED(260, 11),    TO_SIGNED(304, 11),    TO_SIGNED(342, 11),    TO_SIGNED(372, 11),    TO_SIGNED(395, 11),    TO_SIGNED(410, 11),    TO_SIGNED(416, 11),    TO_SIGNED(414, 11),
    TO_SIGNED(403, 11),    TO_SIGNED(384, 11),    TO_SIGNED(358, 11),    TO_SIGNED(325, 11),    TO_SIGNED(285, 11),    TO_SIGNED(240, 11),    TO_SIGNED(190, 11),    TO_SIGNED(137, 11),
    TO_SIGNED(82, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-31, 11),    TO_SIGNED(-86, 11),    TO_SIGNED(-140, 11),    TO_SIGNED(-190, 11),    TO_SIGNED(-235, 11),    TO_SIGNED(-276, 11),
    TO_SIGNED(-311, 11),    TO_SIGNED(-339, 11),    TO_SIGNED(-360, 11),    TO_SIGNED(-374, 11),    TO_SIGNED(-380, 11),    TO_SIGNED(-378, 11),    TO_SIGNED(-368, 11),    TO_SIGNED(-351, 11),
    TO_SIGNED(-328, 11),    TO_SIGNED(-297, 11),    TO_SIGNED(-261, 11),    TO_SIGNED(-220, 11),    TO_SIGNED(-175, 11),    TO_SIGNED(-127, 11),    TO_SIGNED(-77, 11),    TO_SIGNED(-25, 11),
    TO_SIGNED(25, 11),    TO_SIGNED(76, 11),    TO_SIGNED(124, 11),    TO_SIGNED(170, 11),    TO_SIGNED(212, 11),    TO_SIGNED(249, 11),    TO_SIGNED(280, 11),    TO_SIGNED(306, 11),
    TO_SIGNED(325, 11),    TO_SIGNED(338, 11),    TO_SIGNED(343, 11),    TO_SIGNED(342, 11),    TO_SIGNED(334, 11),    TO_SIGNED(318, 11),    TO_SIGNED(297, 11),    TO_SIGNED(270, 11),
    TO_SIGNED(238, 11),    TO_SIGNED(201, 11),    TO_SIGNED(160, 11),    TO_SIGNED(117, 11),    TO_SIGNED(71, 11),    TO_SIGNED(25, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(-66, 11),
    TO_SIGNED(-110, 11),    TO_SIGNED(-151, 11),    TO_SIGNED(-188, 11),    TO_SIGNED(-222, 11),    TO_SIGNED(-250, 11),    TO_SIGNED(-273, 11),    TO_SIGNED(-291, 11),    TO_SIGNED(-302, 11),
    TO_SIGNED(-307, 11),    TO_SIGNED(-306, 11),    TO_SIGNED(-299, 11),    TO_SIGNED(-285, 11),    TO_SIGNED(-266, 11),    TO_SIGNED(-242, 11),    TO_SIGNED(-213, 11),    TO_SIGNED(-181, 11),
    TO_SIGNED(-145, 11),    TO_SIGNED(-106, 11),    TO_SIGNED(-66, 11),    TO_SIGNED(-24, 11),    TO_SIGNED(16, 11),    TO_SIGNED(56, 11),    TO_SIGNED(95, 11),    TO_SIGNED(132, 11),
    TO_SIGNED(165, 11),    TO_SIGNED(195, 11),    TO_SIGNED(220, 11),    TO_SIGNED(241, 11),    TO_SIGNED(256, 11),    TO_SIGNED(266, 11),    TO_SIGNED(271, 11),    TO_SIGNED(270, 11),
    TO_SIGNED(264, 11),    TO_SIGNED(252, 11),    TO_SIGNED(235, 11),    TO_SIGNED(214, 11),    TO_SIGNED(189, 11),    TO_SIGNED(160, 11),    TO_SIGNED(128, 11),    TO_SIGNED(95, 11),
    TO_SIGNED(59, 11),    TO_SIGNED(23, 11),    TO_SIGNED(-12, 11),    TO_SIGNED(-48, 11),    TO_SIGNED(-82, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-143, 11),    TO_SIGNED(-168, 11),
    TO_SIGNED(-191, 11),    TO_SIGNED(-209, 11),    TO_SIGNED(-222, 11),    TO_SIGNED(-231, 11),    TO_SIGNED(-235, 11),    TO_SIGNED(-234, 11),    TO_SIGNED(-229, 11),    TO_SIGNED(-218, 11),
    TO_SIGNED(-204, 11),    TO_SIGNED(-186, 11),    TO_SIGNED(-164, 11),    TO_SIGNED(-139, 11),    TO_SIGNED(-112, 11),    TO_SIGNED(-83, 11),    TO_SIGNED(-52, 11),    TO_SIGNED(-21, 11),
    TO_SIGNED(9, 11),     TO_SIGNED(39, 11),    TO_SIGNED(68, 11),    TO_SIGNED(95, 11),    TO_SIGNED(120, 11),    TO_SIGNED(142, 11),    TO_SIGNED(161, 11),    TO_SIGNED(177, 11),
    TO_SIGNED(188, 11),   TO_SIGNED(195, 11),    TO_SIGNED(199, 11),    TO_SIGNED(198, 11),    TO_SIGNED(193, 11),    TO_SIGNED(185, 11),    TO_SIGNED(173, 11),    TO_SIGNED(157, 11),
    TO_SIGNED(139, 11),   TO_SIGNED(118, 11),    TO_SIGNED(95, 11),    TO_SIGNED(70, 11),    TO_SIGNED(45, 11),    TO_SIGNED(19, 11),    TO_SIGNED(-6, 11),    TO_SIGNED(-31, 11),
    TO_SIGNED(-55, 11),   TO_SIGNED(-78, 11),    TO_SIGNED(-99, 11),    TO_SIGNED(-117, 11),    TO_SIGNED(-132, 11),    TO_SIGNED(-145, 11),    TO_SIGNED(-154, 11),    TO_SIGNED(-160, 11),
    TO_SIGNED(-163, 11),  TO_SIGNED(-162, 11),    TO_SIGNED(-158, 11),    TO_SIGNED(-151, 11),    TO_SIGNED(-141, 11),    TO_SIGNED(-128, 11),    TO_SIGNED(-113, 11),    TO_SIGNED(-96, 11),
    TO_SIGNED(-77, 11),   TO_SIGNED(-58, 11),    TO_SIGNED(-37, 11),    TO_SIGNED(-16, 11),    TO_SIGNED(4, 11),    TO_SIGNED(24, 11),    TO_SIGNED(43, 11),    TO_SIGNED(61, 11),
    TO_SIGNED(77, 11),    TO_SIGNED(91, 11),    TO_SIGNED(104, 11),    TO_SIGNED(113, 11),    TO_SIGNED(120, 11),    TO_SIGNED(125, 11),    TO_SIGNED(127, 11),    TO_SIGNED(126, 11),
    TO_SIGNED(123, 11),   TO_SIGNED(117, 11),    TO_SIGNED(109, 11),    TO_SIGNED(99, 11),    TO_SIGNED(87, 11),    TO_SIGNED(74, 11),    TO_SIGNED(59, 11),    TO_SIGNED(44, 11),
    TO_SIGNED(29, 11),    TO_SIGNED(13, 11),    TO_SIGNED(-2, 11),    TO_SIGNED(-17, 11),    TO_SIGNED(-31, 11),    TO_SIGNED(-44, 11),    TO_SIGNED(-56, 11),    TO_SIGNED(-67, 11),
    TO_SIGNED(-75, 11),   TO_SIGNED(-82, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-90, 11),    TO_SIGNED(-91, 11),    TO_SIGNED(-90, 11),    TO_SIGNED(-87, 11),    TO_SIGNED(-83, 11),
    TO_SIGNED(-77, 11),   TO_SIGNED(-69, 11),    TO_SIGNED(-61, 11),    TO_SIGNED(-51, 11),    TO_SIGNED(-41, 11),    TO_SIGNED(-31, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(-9, 11),
    TO_SIGNED(1, 11),     TO_SIGNED(11, 11),    TO_SIGNED(20, 11),    TO_SIGNED(28, 11),    TO_SIGNED(36, 11),    TO_SIGNED(42, 11),    TO_SIGNED(47, 11),    TO_SIGNED(51, 11),
    TO_SIGNED(54, 11),    TO_SIGNED(55, 11),    TO_SIGNED(55, 11),    TO_SIGNED(54, 11),    TO_SIGNED(51, 11),    TO_SIGNED(48, 11),    TO_SIGNED(44, 11),    TO_SIGNED(39, 11),
    TO_SIGNED(34, 11),    TO_SIGNED(28, 11),    TO_SIGNED(22, 11),    TO_SIGNED(16, 11),    TO_SIGNED(10, 11),    TO_SIGNED(5, 11),    TO_SIGNED(0, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-9, 11),    TO_SIGNED(-13, 11),    TO_SIGNED(-16, 11),    TO_SIGNED(-18, 11),    TO_SIGNED(-19, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(-20, 11),    TO_SIGNED(-20, 11),
    TO_SIGNED(-19, 11),   TO_SIGNED(-18, 11),    TO_SIGNED(-16, 11),    TO_SIGNED(-14, 11),    TO_SIGNED(-11, 11),    TO_SIGNED(-9, 11),    TO_SIGNED(-7, 11),    TO_SIGNED(-5, 11),
    TO_SIGNED(-3, 11),    TO_SIGNED(-2, 11),    TO_SIGNED(0, 11),    TO_SIGNED(0, 11)
  );

  -- QUELQUES PETITES MODIFICATIONS FAITES POUR AIDER VIVADO A FAIRE LES BONS
  -- CHOIX D'IMPLEMENTATION...

  ATTRIBUTE RAM_STYLE : string;
  ATTRIBUTE RAM_STYLE of memory: signal is "BLOCK";

BEGIN

  PROCESS (CLOCK)
  BEGIN
    IF (CLOCK'event AND CLOCK = '1') THEN
      DATA_OUT <= STD_LOGIC_VECTOR( memory(to_integer(UNSIGNED(ADDR_R))) );
    END IF;
  END PROCESS;
  
END Behavioral;